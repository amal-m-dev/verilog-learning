module siso_top (
    si,
    clk,
    rst,
    so);

    
    
endmodule